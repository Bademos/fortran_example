b0VIM 8.2      �j�c)l �  vadique                                 debian                                  ~vadique/homework/lab_3_roma_alloc/src/main.f90                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              utf-8 3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp           ,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ad  t
  @     ,       �  �  �  �  �  �  �  W    �  �  �  �  j  M  (  '  &  %      �  �  �  �  p  6        �  �  �  �  �  �  0    �  �  n  c  _  @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeend program reference_lab_list       ! end if    !   call Output_list(output_file, set3, "Исходный список:", "rewind")       ! call Output_ex(output_file,list, list_comm, "poehali!", "rewind")    ! if (Associated(List1)) then !call Output_list(output_file, List1, "Исходный список:", "rewind")        !call control(set1,set2,set3)  !  end if  !        set3 => set3%next%next  !  if (isContainChar(set3%char, set1,.false.)) then      !  end if  !     call Conjuct(set3,set2)  !  if (.not.isContainChar(set2%char, set1,.false.)) then   ! call setDivide(set1,set2,set3)   ! call setMaking(List2,Set2)  !  call setMaking(List1,Set1)    List2 = Read_list(F2)    List1 = Read_list(F1)        output_file = "output.txt"       input_file  = "../data/input.txt"    F2  = "../data/file2.txt"    F1  = "../data/file1.txt"          Set1,Set2,Set3    type(symbol), allocatable   :: List1, List2,&    logical                   :: isChr    character(kind=CH_)       :: cr = 'u'    integer                   :: num_bracket = 0,pos = 1    character(:), allocatable :: input_file, output_file, F1, F2, F4    implicit none     use List_IO    use  List_Process    use Environment program reference_lab_list  